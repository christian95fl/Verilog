module inv (input A, output B);
wire A;
wire B;
  assign B = ~A;
endmodule //
