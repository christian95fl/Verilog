module fport(output [3:0] data);
  wire [3:0] data;
  assign data = 4'b1010;
endmodule //
