`difine F_1Hz 12_000_000
